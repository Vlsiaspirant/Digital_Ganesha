
`timescale 1ns / 1ps

module ganesha(
    input wire clk,en,
    input [4:0]address,
    output reg [63:0]data_out
    );
    
    reg [63:0]register[31:0];
    initial begin 
    data_out = 64'd0;
    end 
    
    initial begin 
    
        register[0]  = 64'b0000000000000000000000000000000000000000000000000000000000000000;
        register[1]  = 64'b0000000000000000000000000000000000000000000000000000000000000000;
        register[2]  = 64'b0000000000000000000000000000000000000000000000000000000000000000; 
        register[3]  = 64'b0000000000000000000000000000000000000000000000000000000000000000;
        register[4]  = 64'b0000000000000000000000100100000000000000000000000000000000001111;
        register[5]  = 64'b0000000000000000000001110100000000000000000000000000000000001111;
        register[6]  = 64'b0000000000000000000011111100000000000000000000011111110000001111; 
        register[7]  = 64'b0000000000000000000001110100001111111111111000100000001000001111;
        register[8]  = 64'b0001111111111110000000100100010000000000000100100000000100001111;
        register[9]  = 64'b0010000000000001000000000100100000000000000010010000000100001111;
       register[10] = 64'b0100000000000010000011111101000000000000000001010000000010001111; 
       register[11] = 64'b0010000000000100000100000010000000000000000000110000000010001111;
       register[12] = 64'b0001000000001000001000000010000000000000000000010000000010001111;
       register[13] = 64'b0000111111111000010000000000000000000000000000010000000010001111;
       register[14] = 64'b0001000000000100100000000000000000000000000000010000000010001111;
       register[15] = 64'b0011000000000010100000000000001100000000000000010000000001111111; 
       register[16] = 64'b0111000100000001000000000000000010000000000000010000000000111111;
       register[17] = 64'b1111000000000000111111111111111100000000000000010000000000011111;
       register[18] = 64'b0111000100000001000000000000000000000000000000010000000111101111;
       register[19] = 64'b0011000000000010100000000000000000000000000000010000001000001111; 
       register[20] = 64'b0001000000000100010000000000000000000000000000010000000100001111;
       register[21] = 64'b0000111111111000001000000010000000000000000000010000000010001111;
       register[22] = 64'b0001000000001000000100000010000000000000000000110000000010001111;
       register[23] = 64'b0010000000000100000001111101000000000000000001010000000010001111; 
       register[24] = 64'b0100000000000010000000000010100000000000000010010000000010001111;
       register[25] = 64'b0100000000000001000000111110010000000000000100100000000010001111;
       register[26] = 64'b0011111111111110000000111110001111111111111001000000000100001111;
       register[27] = 64'b0000000000000000000000000010000000000000000000100000000100001111; 
       register[28] = 64'b0000000000000000000000000000000000000000000000100000001000001111;
       register[29] = 64'b0000000000000000000000000000000000000000000000011111110000001111;
       register[30] = 64'b0000000000000000000000000000000000000000000000000000000000001111;
       register[31] = 64'b0000000000000000000000000000000000000000000000000000000100001111; 
    end 
    
    always @ (posedge clk) begin 
    
    if (en==1'b1)
     data_out <= register[address];  
     else 
     data_out <= 64'd0;
    end
    
endmodule
